`timescale 1ns/1ns

module dds_tb();
    logic clk, rst;
    logic [7:0] out;
    dds dd(clk, rst, out);
    initial begin
		clk = 0;
		forever #5 clk = ~clk;
	end

    initial begin
        rst = 1;
        #5;
        rst = 0;

	#3000;
	#100 $stop;
    end

endmodule