`timescale 1ns/1ns

module messageprocess_tb();
    logic clk, rst, send;
    logic [4:0] msg;
    logic SerOut;
    messageProcess_TOP messageProcess_TOP(clk, rst, send, msg,  SerOut);
    initial begin
		clk = 0;
		forever #5 clk = ~clk;
	end

    initial begin
        rst = 1;
        msg = 5'b10110;
        send = 0;
        #7;
        rst = 0;
        #10
        send = 1;

        #10
        send = 0;


	#1000000 $stop;
    end

endmodule