module zero(output out);

	assign out = 0;


endmodule

module one(output out);

	assign out = 1;


endmodule

module m128(output [7:0]out);
	assign out = 8'd128;

endmodule

